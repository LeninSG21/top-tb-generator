module ALU #(parameter W = 9, parameter H = 2'h12)(
    input x, output y, input [3:0] zz, output[W-1:0]yy);